module incr2();



endmodule