module opDecode(instruct);
	input [15:0] instruct;
	



endmodule